`timescale 1ns / 1ps
module CPU(
input CLK100MHZ

);


CONTROL_UNIT CU_I(




);






endmodule
